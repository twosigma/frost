/*
 *    Copyright 2026 Two Sigma Open Source, LLC
 *
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *
 *        http://www.apache.org/licenses/LICENSE-2.0
 *
 *    Unless required by applicable law or agreed to in writing, software
 *    distributed under the License is distributed on an "AS IS" BASIS,
 *    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *    See the License for the specific language governing permissions and
 *    limitations under the License.
 */

/*
  Instruction Decode (ID) stage - Third stage of the 6-stage RISC-V pipeline.
  This module decodes RISC-V instructions into control signals and immediate values.
  It instantiates decoders for instruction type determination and immediate
  value extraction. The module identifies load instructions, store operations, branch
  conditions, and ALU operations. It supports pipeline flushing on branch mispredictions
  and stalling for hazards. The decoded information is passed to the Execute stage through
  a pipeline register that can be flushed or stalled as needed for correct program execution.
*/
module id_stage #(
    parameter int unsigned XLEN = 32
) (
    input logic i_clk,
    input riscv_pkg::pipeline_ctrl_t i_pipeline_ctrl,
    input riscv_pkg::from_pd_to_id_t i_from_pd_to_id,
    input riscv_pkg::rf_to_fwd_t i_rf_to_id,  // Regfile read data (combinational from PD src regs)
    input riscv_pkg::from_ma_to_wb_t i_from_ma_to_wb,  // WB bypass (WB writes same cycle ID reads)
    output riscv_pkg::from_id_to_ex_t o_from_id_to_ex
);

  // Internal signals for decoded instruction information
  riscv_pkg::instr_t instruction;
  riscv_pkg::instr_op_e instruction_operation;
  riscv_pkg::branch_taken_op_e branch_operation;
  riscv_pkg::store_op_e store_operation;
  logic is_load_instruction;
  // Immediate values for different instruction formats
  logic [31:0] immediate_i_type;  // I-type immediate
  logic [31:0] immediate_s_type;  // S-type immediate (for stores)
  logic [31:0] immediate_b_type;  // B-type immediate (for branches)
  logic [31:0] immediate_u_type;  // U-type immediate (upper 20 bits)
  logic [31:0] immediate_j_type;  // J-type immediate (for jumps)

  assign instruction = i_from_pd_to_id.instruction;

  // Instantiate instruction decoder to determine operation type
  instr_decoder instr_decoder_inst (
      .i_instr(instruction),
      .o_instr_op(instruction_operation),
      .o_store_op(store_operation),
      .o_branch_taken_op(branch_operation)
  );

  // Extract and sign-extend immediate values from instruction fields
  // I-type: 12-bit immediate in bits [31:20]
  assign immediate_i_type = {
    {20{instruction.funct7[6]}}, instruction.funct7, instruction.source_reg_2
  };
  // S-type: 12-bit immediate split between bits [31:25] and [11:7]
  assign immediate_s_type = {{20{instruction.funct7[6]}}, instruction.funct7, instruction.dest_reg};
  // B-type: 13-bit immediate (branch offset) scrambled in instruction
  assign immediate_b_type = {
    {19{instruction.funct7[6]}},
    instruction.funct7[6],
    instruction.dest_reg[0],
    instruction.funct7[5:0],
    instruction.dest_reg[4:1],
    1'b0
  };
  // U-type: 20-bit immediate in upper bits, lower 12 bits are zero
  assign immediate_u_type = {instruction[31:12], 12'h0};
  // J-type: 21-bit jump offset scrambled in instruction
  assign immediate_j_type = {
    {11{instruction[31]}},
    instruction[31],
    instruction[19:12],
    instruction[20],
    instruction[30:21],
    1'b0
  };

  assign is_load_instruction = instruction.opcode == riscv_pkg::OPC_LOAD;

  // Direct decode of load type from instruction bits (parallel with instruction_operation)
  // This breaks the dependency chain: instruction → instruction_operation → is_load_*
  // Load funct3: 000=LB, 001=LH, 010=LW, 100=LBU, 101=LHU
  logic is_load_byte_direct;
  logic is_load_halfword_direct;
  logic is_load_unsigned_direct;
  assign is_load_byte_direct = is_load_instruction &&
                               (instruction.funct3 == 3'b000 || instruction.funct3 == 3'b100);
  assign is_load_halfword_direct = is_load_instruction &&
                                   (instruction.funct3 == 3'b001 || instruction.funct3 == 3'b101);
  assign is_load_unsigned_direct = is_load_instruction && instruction.funct3[2];

  // Direct decode of multiply/divide from instruction bits
  // M-extension uses opcode=OP (0110011), funct7=0000001
  logic is_m_extension;
  logic is_multiply_direct;
  logic is_divide_direct;
  assign is_m_extension = (instruction.opcode == riscv_pkg::OPC_OP) &&
                          (instruction.funct7 == 7'b0000001);
  assign is_multiply_direct = is_m_extension && !instruction.funct3[2];  // funct3[2]=0 for MUL*
  assign is_divide_direct = is_m_extension && instruction.funct3[2];  // funct3[2]=1 for DIV/REM

  // CSR instruction detection and field extraction (Zicsr extension)
  logic is_csr_instruction;
  logic [11:0] csr_address;
  logic [4:0] csr_imm;
  assign is_csr_instruction = instruction.opcode == riscv_pkg::OPC_CSR;
  assign csr_address = {
    instruction.funct7, instruction.source_reg_2
  };  // CSR address in bits [31:20]
  assign csr_imm = instruction.source_reg_1;  // Zero-extended immediate for CSRRWI/CSRRSI/CSRRCI

  // A extension (atomics) detection - decode directly from instruction bits
  logic is_amo_instruction;
  logic is_lr;
  logic is_sc;
  assign is_amo_instruction = instruction.opcode == riscv_pkg::OPC_AMO;
  // LR.W: funct7[6:2]=00010, funct3=010
  // SC.W: funct7[6:2]=00011, funct3=010
  assign is_lr = is_amo_instruction && (instruction.funct3 == 3'b010) &&
                 (instruction.funct7[6:2] == 5'b00010);
  assign is_sc = is_amo_instruction && (instruction.funct3 == 3'b010) &&
                 (instruction.funct7[6:2] == 5'b00011);

  // Privileged instruction detection - decode directly from instruction bits
  // All use opcode=SYSTEM (1110011), funct3=000
  logic is_mret;
  logic is_wfi;
  logic is_ecall;
  logic is_ebreak;
  logic is_priv_instruction;
  assign is_priv_instruction = (instruction.opcode == riscv_pkg::OPC_CSR) &&
                               (instruction.funct3 == 3'b000);
  // ECALL: funct7=0000000, rs2=00000
  assign is_ecall = is_priv_instruction &&
                    (instruction.funct7 == 7'b0000000) && (instruction.source_reg_2 == 5'b00000);
  // EBREAK: funct7=0000000, rs2=00001
  assign is_ebreak = is_priv_instruction &&
                     (instruction.funct7 == 7'b0000000) && (instruction.source_reg_2 == 5'b00001);
  // MRET: funct7=0011000, rs2=00010
  assign is_mret = is_priv_instruction &&
                   (instruction.funct7 == 7'b0011000) && (instruction.source_reg_2 == 5'b00010);
  // WFI: funct7=0001000, rs2=00101
  assign is_wfi = is_priv_instruction &&
                  (instruction.funct7 == 7'b0001000) && (instruction.source_reg_2 == 5'b00101);

  // Direct decode of JAL/JALR for timing - don't depend on instruction_operation
  logic is_jal_direct;
  logic is_jalr_direct;
  assign is_jal_direct = instruction.opcode == riscv_pkg::OPC_JAL;
  assign is_jalr_direct = (instruction.opcode == riscv_pkg::OPC_JALR) &&
                          (instruction.funct3 == 3'b000);

  // ===========================================================================
  // TIMING OPTIMIZATION: Pre-compute RAS instruction type detection
  // ===========================================================================
  // These flags are computed here (ID stage) from registered inputs and passed
  // to EX stage to remove comparisons from the critical ras_correct path.
  //
  // is_ras_return: JALR with rs1 in {x1, x5}, rd = x0, imm = 0
  // is_ras_call: JAL/JALR with rd in {x1, x5}
  // ras_predicted_target_nonzero: ras_predicted_target != 0

  logic is_ras_return_precomputed;
  logic is_ras_call_precomputed;
  logic rs1_is_link_reg;
  logic rd_is_link_reg;

  assign rs1_is_link_reg = (instruction.source_reg_1 == 5'd1) || (instruction.source_reg_1 == 5'd5);
  assign rd_is_link_reg = (instruction.dest_reg == 5'd1) || (instruction.dest_reg == 5'd5);

  // Return: JALR with rs1 in {x1, x5}, rd = x0, imm = 0
  // The immediate for JALR is in I-type format: funct7[6:0] ++ source_reg_2[4:0]
  assign is_ras_return_precomputed = is_jalr_direct &&
                                     rs1_is_link_reg &&
                                     (instruction.dest_reg == 5'd0) &&
                                     (immediate_i_type == 32'b0);

  // Call: JAL or JALR with rd in {x1, x5}
  assign is_ras_call_precomputed = (is_jal_direct || is_jalr_direct) && rd_is_link_reg;

  // TIMING OPTIMIZATION: Pre-compute expected rs1 for RAS target verification.
  // For JALR returns: actual_target = rs1 + immediate_i_type
  // Therefore: expected_rs1 = ras_predicted_target - immediate_i_type
  // This allows EX stage to verify RAS prediction by comparing forwarded_rs1
  // with this pre-computed value, removing the JALR adder from the critical path.
  logic [XLEN-1:0] ras_expected_rs1_precomputed;
  assign ras_expected_rs1_precomputed = i_from_pd_to_id.ras_predicted_target -
                                        XLEN'(signed'(immediate_i_type));

  // ===========================================================================
  // TIMING OPTIMIZATION: Pre-compute BTB target verification
  // ===========================================================================
  // Same algebraic transformation as RAS, applied to BTB comparison.
  // For JALR: btb_expected_rs1 = btb_predicted_target - immediate_i_type
  //   EX stage compares: forwarded_rs1 == btb_expected_rs1
  // For non-JALR (JAL/branches): targets are PC-relative, computed here
  //   Compare precomputed target with btb_predicted_target in ID stage
  //   This removes the entire comparison from EX stage critical path
  logic [XLEN-1:0] btb_expected_rs1_precomputed;
  assign btb_expected_rs1_precomputed = i_from_pd_to_id.btb_predicted_target -
                                        XLEN'(signed'(immediate_i_type));

  // For non-JALR, select the appropriate precomputed target
  // JAL uses jal_target_precomputed, branches use branch_target_precomputed
  logic [XLEN-1:0] precomputed_target_for_btb;
  assign precomputed_target_for_btb = is_jal_direct ?
                                      jal_target_precomputed : branch_target_precomputed;

  // Pre-compute BTB correctness for non-JALR instructions
  // This comparison happens in ID stage where timing is not critical
  logic btb_correct_non_jalr_precomputed;
  assign btb_correct_non_jalr_precomputed = (precomputed_target_for_btb ==
                                             i_from_pd_to_id.btb_predicted_target);

  // Pre-computed branch/jump targets for pipeline balancing.
  // Computing PC-relative targets here removes adders from EX stage critical path.
  // Only JALR target is computed in EX since it requires forwarded rs1.
  logic [XLEN-1:0] branch_target_precomputed;
  logic [XLEN-1:0] jal_target_precomputed;
  assign branch_target_precomputed = i_from_pd_to_id.program_counter +
                                     XLEN'(signed'(immediate_b_type));
  assign jal_target_precomputed = i_from_pd_to_id.program_counter +
                                  XLEN'(signed'(immediate_j_type));

  // WB bypass for regfile data: When WB writes to a register that ID is reading,
  // we must use the WB write data instead of the regfile read data. This is because
  // the regfile read (async) happens the same cycle as the WB write (sync), so the
  // regfile read would get stale data before the write commits.
  logic wb_bypass_rs1;
  logic wb_bypass_rs2;
  logic [XLEN-1:0] source_reg_1_data_bypassed;
  logic [XLEN-1:0] source_reg_2_data_bypassed;

  assign wb_bypass_rs1 = i_from_ma_to_wb.regfile_write_enable &&
                         |i_from_ma_to_wb.instruction.dest_reg &&
                         (i_from_ma_to_wb.instruction.dest_reg ==
                          i_from_pd_to_id.source_reg_1_early);
  assign wb_bypass_rs2 = i_from_ma_to_wb.regfile_write_enable &&
                         |i_from_ma_to_wb.instruction.dest_reg &&
                         (i_from_ma_to_wb.instruction.dest_reg ==
                          i_from_pd_to_id.source_reg_2_early);

  assign source_reg_1_data_bypassed = wb_bypass_rs1 ? i_from_ma_to_wb.regfile_write_data :
                                                      i_rf_to_id.source_reg_1_data;
  assign source_reg_2_data_bypassed = wb_bypass_rs2 ? i_from_ma_to_wb.regfile_write_data :
                                                      i_rf_to_id.source_reg_2_data;

  // TIMING OPTIMIZATION: Pre-compute x0 check for source registers.
  // This moves the ~|source_reg NOR gate out of the EX stage critical path.
  // The forwarding unit uses these registered flags instead of computing them combinationally.
  logic source_reg_1_is_x0;
  logic source_reg_2_is_x0;
  assign source_reg_1_is_x0 = ~|i_from_pd_to_id.source_reg_1_early;
  assign source_reg_2_is_x0 = ~|i_from_pd_to_id.source_reg_2_early;

  // Pipeline register: latch decoded values and pass to Execute stage
  always_ff @(posedge i_clk) begin
    // On reset, insert a NOP (no operation) into the pipeline
    if (i_pipeline_ctrl.reset) begin
      o_from_id_to_ex.instruction                  <= riscv_pkg::NOP;
      o_from_id_to_ex.instruction_operation        <= riscv_pkg::ADDI;  // ADDI x0, x0, 0 (NOP)
      o_from_id_to_ex.is_load_instruction          <= 1'b0;
      o_from_id_to_ex.is_load_byte                 <= 1'b0;
      o_from_id_to_ex.is_load_halfword             <= 1'b0;
      o_from_id_to_ex.is_load_unsigned             <= 1'b0;
      o_from_id_to_ex.is_multiply                  <= 1'b0;
      o_from_id_to_ex.is_divide                    <= 1'b0;
      o_from_id_to_ex.program_counter              <= '0;
      o_from_id_to_ex.branch_operation             <= riscv_pkg::NULL;
      o_from_id_to_ex.store_operation              <= riscv_pkg::STN;  // Store nothing
      o_from_id_to_ex.is_jump_and_link             <= 1'b0;
      o_from_id_to_ex.is_jump_and_link_register    <= 1'b0;
      o_from_id_to_ex.is_csr_instruction           <= 1'b0;
      o_from_id_to_ex.csr_address                  <= '0;
      o_from_id_to_ex.csr_imm                      <= '0;
      // A extension (atomics)
      o_from_id_to_ex.is_amo_instruction           <= 1'b0;
      o_from_id_to_ex.is_lr                        <= 1'b0;
      o_from_id_to_ex.is_sc                        <= 1'b0;
      // Privileged instructions (trap handling)
      o_from_id_to_ex.is_mret                      <= 1'b0;
      o_from_id_to_ex.is_wfi                       <= 1'b0;
      o_from_id_to_ex.is_ecall                     <= 1'b0;
      o_from_id_to_ex.is_ebreak                    <= 1'b0;
      o_from_id_to_ex.link_address                 <= '0;
      // Pre-computed branch/jump targets (pipeline balancing)
      o_from_id_to_ex.branch_target_precomputed    <= '0;
      o_from_id_to_ex.jal_target_precomputed       <= '0;
      // Regfile read data (read in ID stage using early source regs from PD)
      o_from_id_to_ex.source_reg_1_data            <= '0;
      o_from_id_to_ex.source_reg_2_data            <= '0;
      // Pre-computed x0 check flags (timing optimization)
      o_from_id_to_ex.source_reg_1_is_x0           <= 1'b1;  // NOP uses x0
      o_from_id_to_ex.source_reg_2_is_x0           <= 1'b1;  // NOP uses x0
      // Branch prediction metadata
      o_from_id_to_ex.btb_hit                      <= 1'b0;
      o_from_id_to_ex.btb_predicted_taken          <= 1'b0;
      o_from_id_to_ex.btb_predicted_target         <= '0;
      // RAS prediction metadata
      o_from_id_to_ex.ras_predicted                <= 1'b0;
      o_from_id_to_ex.ras_predicted_target         <= '0;
      o_from_id_to_ex.ras_checkpoint_tos           <= '0;
      o_from_id_to_ex.ras_checkpoint_valid_count   <= '0;
      // TIMING OPTIMIZATION: Pre-computed RAS instruction type flags
      o_from_id_to_ex.is_ras_return                <= 1'b0;
      o_from_id_to_ex.is_ras_call                  <= 1'b0;
      o_from_id_to_ex.ras_predicted_target_nonzero <= 1'b0;
      o_from_id_to_ex.ras_expected_rs1             <= '0;
      // TIMING OPTIMIZATION: Pre-computed BTB verification
      o_from_id_to_ex.btb_correct_non_jalr         <= 1'b0;
      o_from_id_to_ex.btb_expected_rs1             <= '0;
    end else if (~i_pipeline_ctrl.stall) begin
      // When pipeline is not stalled, pass decoded instruction to Execute stage
      // If flushing (e.g., due to branch), insert NOP instead
      o_from_id_to_ex.instruction <= i_pipeline_ctrl.flush ? riscv_pkg::NOP : instruction;
      o_from_id_to_ex.instruction_operation <= i_pipeline_ctrl.flush ? riscv_pkg::ADDI :
                                                                       instruction_operation;
      o_from_id_to_ex.is_load_instruction <= i_pipeline_ctrl.flush ? 1'b0 : is_load_instruction;
      // Determine load size and sign extension - use direct decode for timing
      o_from_id_to_ex.is_load_byte <= i_pipeline_ctrl.flush ? 1'b0 : is_load_byte_direct;
      o_from_id_to_ex.is_load_halfword <= i_pipeline_ctrl.flush ? 1'b0 : is_load_halfword_direct;
      o_from_id_to_ex.is_load_unsigned <= i_pipeline_ctrl.flush ? 1'b0 : is_load_unsigned_direct;
      // Check if this is a multiply operation (M extension) - use direct decode
      o_from_id_to_ex.is_multiply <= i_pipeline_ctrl.flush ? 1'b0 : is_multiply_direct;
      // Check if this is a divide/remainder operation (M extension) - use direct decode
      o_from_id_to_ex.is_divide <= i_pipeline_ctrl.flush ? 1'b0 : is_divide_direct;
      o_from_id_to_ex.program_counter <= i_from_pd_to_id.program_counter;
      o_from_id_to_ex.branch_operation <= i_pipeline_ctrl.flush ? riscv_pkg::NULL :
                                                                  branch_operation;
      o_from_id_to_ex.store_operation <= i_pipeline_ctrl.flush ? riscv_pkg::STN : store_operation;
      o_from_id_to_ex.is_jump_and_link <= i_pipeline_ctrl.flush ? 1'b0 : is_jal_direct;
      o_from_id_to_ex.is_jump_and_link_register <= i_pipeline_ctrl.flush ? 1'b0 : is_jalr_direct;
      // CSR instruction fields (Zicsr extension)
      o_from_id_to_ex.is_csr_instruction <= i_pipeline_ctrl.flush ? 1'b0 : is_csr_instruction;
      o_from_id_to_ex.csr_address <= csr_address;
      o_from_id_to_ex.csr_imm <= csr_imm;
      // A extension (atomics)
      o_from_id_to_ex.is_amo_instruction <= i_pipeline_ctrl.flush ? 1'b0 : is_amo_instruction;
      o_from_id_to_ex.is_lr <= i_pipeline_ctrl.flush ? 1'b0 : is_lr;
      o_from_id_to_ex.is_sc <= i_pipeline_ctrl.flush ? 1'b0 : is_sc;
      // Privileged instructions (trap handling)
      o_from_id_to_ex.is_mret <= i_pipeline_ctrl.flush ? 1'b0 : is_mret;
      o_from_id_to_ex.is_wfi <= i_pipeline_ctrl.flush ? 1'b0 : is_wfi;
      o_from_id_to_ex.is_ecall <= i_pipeline_ctrl.flush ? 1'b0 : is_ecall;
      o_from_id_to_ex.is_ebreak <= i_pipeline_ctrl.flush ? 1'b0 : is_ebreak;
      // Pre-computed link address from IF stage
      o_from_id_to_ex.link_address <= i_from_pd_to_id.link_address;
      // Pre-computed branch/jump targets (computed here, used by EX stage)
      o_from_id_to_ex.branch_target_precomputed <= branch_target_precomputed;
      o_from_id_to_ex.jal_target_precomputed <= jal_target_precomputed;
      // Branch prediction metadata - clear on flush (prediction for flushed instr is invalid)
      o_from_id_to_ex.btb_hit <= i_pipeline_ctrl.flush ? 1'b0 : i_from_pd_to_id.btb_hit;
      o_from_id_to_ex.btb_predicted_taken <= i_pipeline_ctrl.flush ? 1'b0 :
                                              i_from_pd_to_id.btb_predicted_taken;
      o_from_id_to_ex.btb_predicted_target <= i_from_pd_to_id.btb_predicted_target;
      // RAS prediction metadata - clear on flush (prediction for flushed instr is invalid)
      o_from_id_to_ex.ras_predicted <= i_pipeline_ctrl.flush ? 1'b0 : i_from_pd_to_id.ras_predicted;
      o_from_id_to_ex.ras_predicted_target <= i_from_pd_to_id.ras_predicted_target;
      o_from_id_to_ex.ras_checkpoint_tos <= i_from_pd_to_id.ras_checkpoint_tos;
      o_from_id_to_ex.ras_checkpoint_valid_count <= i_from_pd_to_id.ras_checkpoint_valid_count;
      // TIMING OPTIMIZATION: Pre-computed RAS instruction type flags
      // These remove comparisons from the EX stage critical path
      o_from_id_to_ex.is_ras_return <= i_pipeline_ctrl.flush ? 1'b0 : is_ras_return_precomputed;
      o_from_id_to_ex.is_ras_call <= i_pipeline_ctrl.flush ? 1'b0 : is_ras_call_precomputed;
      o_from_id_to_ex.ras_predicted_target_nonzero <= |i_from_pd_to_id.ras_predicted_target;
      // Pre-computed expected rs1 for RAS verification (removes JALR adder from critical path)
      o_from_id_to_ex.ras_expected_rs1 <= ras_expected_rs1_precomputed;
      // TIMING OPTIMIZATION: Pre-computed BTB verification
      // For non-JALR: target comparison done in ID stage (no forwarding dependency)
      // For JALR: use btb_expected_rs1 in EX stage (same algebraic transformation as RAS)
      o_from_id_to_ex.btb_correct_non_jalr <= i_pipeline_ctrl.flush ? 1'b0 :
                                              btb_correct_non_jalr_precomputed;
      o_from_id_to_ex.btb_expected_rs1 <= btb_expected_rs1_precomputed;
    end
    // Pass immediate values and regfile data (datapath, not affected by reset - only by stall)
    if (~i_pipeline_ctrl.stall) begin
      o_from_id_to_ex.immediate_u_type   <= immediate_u_type;
      o_from_id_to_ex.immediate_s_type   <= immediate_s_type;
      o_from_id_to_ex.immediate_i_type   <= immediate_i_type;
      o_from_id_to_ex.immediate_b_type   <= immediate_b_type;
      o_from_id_to_ex.immediate_j_type   <= immediate_j_type;
      // Regfile read data (read in ID stage, with WB bypass, registered here for EX stage)
      o_from_id_to_ex.source_reg_1_data  <= source_reg_1_data_bypassed;
      o_from_id_to_ex.source_reg_2_data  <= source_reg_2_data_bypassed;
      // Pre-computed x0 check flags (timing optimization for forwarding unit)
      o_from_id_to_ex.source_reg_1_is_x0 <= source_reg_1_is_x0;
      o_from_id_to_ex.source_reg_2_is_x0 <= source_reg_2_is_x0;
    end
  end

endmodule : id_stage
